module DisplayUnit(clk, lcd_e, lcd_rs, lcd_rw, reset, cs1, cs2, lcd_data,,G_SENSOR_CS_N,G_SENSOR_INT,I2C_SCLK,I2C_SDAT,KEY);

	input G_SENSOR_INT;
	input [1:0]KEY;
	output wire G_SENSOR_CS_N,I2C_SCLK;
	inout I2C_SDAT;
	wire [7:0] LED;
	
	input clk;

	output reg lcd_e, lcd_rs, lcd_rw;
	output reg cs1, cs2, reset;
	output reg [7:0]lcd_data;
	
	//parameter k=18;
	reg [60:0]divider;
	reg [8:0] count;
	reg already_on=0;
	reg[7:0] mem[0:7][0:255];
	reg[7:0] temp1, temp2, temp3, temp4, temp5, temp6, temp7;

	//Raaz variables 
	reg[7:0] tmem[0:7][0:127]; //temporary memory for gameover and welcome
	reg gameover=0; 
	integer l,j, k; 
	reg[7:0] temp_t; 
	integer move_t=0; 
	reg clk_1, clk_2, clk_3, clk_4, clk_5, clk_6, clk_7; 
	integer level=0; 
	integer i1, j1; 
	reg init_w=0, init_g=1; // if init is low that part is executed : w for WELCOME, g for GAMEOVER
	reg start=1; 
	reg [7:0]carmem [8][6]; 
	reg [2:0]car_page=3; 
	integer rate=1; 
	integer ic, jc; 
	wire [1:0]speed;
	integer timer1=0;

	//Pendi's variables
	integer move1=0, move2 =0 , move3 = 0, move4= 0, move5 =0, move6 = 0, move7 = 0;
	integer timer = 0 ;
	integer init1 = 0, init2 =0 ,init3 =0, init4 = 0, init5 =0, init6 = 0, init7 = 0;
	integer col = 0;
	integer i = 0;
	integer page = 0;

DE0_NANO_G_Sensor Sensor(clk,LED,KEY,G_SENSOR_CS_N,G_SENSOR_INT,I2C_SCLK,I2C_SDAT );	
		
//Level update
always@(*) begin
start = (timer1<=50) ? 1 :0 ; 
if(timer<=200) level<=0; 
else if(timer >200 && timer<=500) level<=1; 
else if(timer >5000) level<=2; 
else if(timer >750) level<=3;

clk_1<=divider[22-level] ; 
clk_2<=divider[20-level] ; 
clk_3<=divider[22-level] ; 
clk_4<=divider[22-level] ; 
clk_5<=divider[22-level] ; 
clk_6<=divider[20-level] ; 
clk_7<=divider[22-level] ; 

end

//G Sensor LED Output	
always @(LED) begin 
 if(LED[7]) car_page = 7; 
 else if(LED[6]) car_page = 6;
 else if(LED[5]) car_page = 5;
 else if( (LED [4]) | (LED [3])) car_page = 4;
 else if (LED [2]) car_page = 3 ;
 else if (LED [1]) car_page = 2 ;
 else if (LED [0]) car_page = 1 ; 
 end



// Removed this line assign speed = (rate>0)? rate : -1*rate ; 

//Car Memory Update 
always@(divider[40])begin
	/*if (rate<0 && car_page>=2)car_page =car_page-1; 
	else if (rate>0 && car_page<=7)car_page=car_page+1; */
	for (ic=0; ic<=7; ic=ic+1) begin 
		for (jc=0; jc<=5; jc=jc+1) begin 
			carmem[ic][jc]=0;
		end 
	end
	carmem[car_page][0][5:0]=33; 
	carmem[car_page][1][5:0]=63; 
	carmem[car_page][2][5:0]=63; 
	carmem[car_page][3][5:0]=63; 
	carmem[car_page][4][5:0]=30; 
	carmem[car_page][5][5:0]=12; 
	end
	
// WORD SCORE
	always@(*) begin
	//Clock Symbol -- Score lettering should come here..
	
	//Letter "S"
	mem[0][55][4:0] = 5'b10010; 
	mem[0][56][4:0] = 5'b10101; 
	mem[0][57][4:0] = 5'b10101; 
	mem[0][58][4:0] = 5'b10101; 
	mem[0][59][4:0] = 5'b01001;

	//Letter "C"
	mem[0][61][4:0] = 5'b00100; 
	mem[0][62][4:0] = 5'b01010; 
	mem[0][63][4:0] = 5'b10001;
	mem[0][64][4:0] = 5'b10001;
	mem[0][65][4:0] = 5'b10001;
	
	//Letter "O"
	mem[0][67][4:0] = 5'b01110; 
	mem[0][68][4:0] = 5'b10001; 
	mem[0][69][4:0] = 5'b10001;
	mem[0][70][4:0] = 5'b10001;
	mem[0][71][4:0] = 5'b01110;
	
	//Letter "R"
	mem[0][73][4:0] = 5'b11111; 
	mem[0][74][4:0] = 5'b00101; 
	mem[0][75][4:0] = 5'b00101;
	mem[0][76][4:0] = 5'b01010;
	mem[0][77][4:0] = 5'b10000;
	
	//Letter "E"
	mem[0][79][4:0] = 5'b11111; 
	mem[0][80][4:0] = 5'b10101; 
	mem[0][81][4:0] = 5'b10101;
	mem[0][82][4:0] = 5'b10101;
	mem[0][83][4:0] = 5'b10001;

	
	
	//Colon
	mem[0][85][4:0] = 5'b01010;
	
	for(l=0; l<=127 ; l=l+1) begin 
	tmem[0][l][4:0] = mem [0][l][4:0]; 
	end
	end


	
//Score increasing block			Change in divider[**] ** accordingly for rate of increase of score
	always@(negedge divider[20]) begin //timer 1 to start the process !!!!!
	timer1 = (timer1 >70)? 71 : timer1+1; 
	timer = (timer1<50|timer == 999999)? 0 : (timer +1) ;
	//gameover = (timer>=500)? 1 : 0 ;  
	//Timer digit 100,000's
	if(!gameover)
	begin 
		case(timer/100000)
	0:
		begin
		mem[0][100][4:0] = 5'b01110;
		mem[0][99][4:0] = 5'b10001;
		mem[0][98][4:0] = 5'b10001;
		mem[0][97][4:0] = 5'b01110;
		end
	1:
		begin
		mem[0][100][4:0] = 5'b10000;
		mem[0][99][4:0] = 5'b11111;
		mem[0][98][4:0] = 5'b10010;
		mem[0][97][4:0] = 5'b00000;
		end
	2:
		begin
		mem[0][100][4:0] = 5'b10010;
		mem[0][99][4:0] = 5'b10101;
		mem[0][98][4:0] = 5'b11001;
		mem[0][97][4:0] = 5'b10010;
		end
	3:
		begin
		mem[0][100][4:0] = 5'b01010;
		mem[0][99][4:0] = 5'b10101;
		mem[0][98][4:0] = 5'b10101;
		mem[0][97][4:0] = 5'b10001;		
		end
	4:
	begin
		mem[0][100][4:0] = 5'b11111;
		mem[0][99][4:0] = 5'b01010;
		mem[0][98][4:0] = 5'b01100;
		mem[0][97][4:0] = 5'b01000;	
	end
	5:
	begin
		mem[0][100][4:0] = 5'b01001;
		mem[0][99][4:0] = 5'b10101;
		mem[0][98][4:0] = 5'b10101;
		mem[0][97][4:0] = 5'b10111;
	end
	6:
	begin
		mem[0][100][4:0] = 5'b01000;
		mem[0][99][4:0] = 5'b10101;
		mem[0][98][4:0] = 5'b10101;
		mem[0][97][4:0] = 5'b01110;
	end
	7:
	begin
		mem[0][100][4:0] = 5'b00011;
		mem[0][99][4:0] = 5'b00101;
		mem[0][98][4:0] = 5'b01001;
		mem[0][97][4:0] = 5'b10001;
	end
	
	8:
	begin
		mem[0][100][4:0] = 5'b01010;
		mem[0][99][4:0] = 5'b10101;
		mem[0][98][4:0] = 5'b10101;
		mem[0][97][4:0] = 5'b01010;
	end
	9: begin
		mem[0][100][4:0] = 5'b01110;
		mem[0][99][4:0] = 5'b10101;
		mem[0][98][4:0] = 5'b10101;
		mem[0][97][4:0] = 5'b00010;
		end
	default : 
		begin
		mem[0][100][4:0] = 5'b01110;
		mem[0][99][4:0] = 5'b10001;
		mem[0][98][4:0] = 5'b10001;
		mem[0][97][4:0] = 5'b01110;
	end
	endcase
	
	
	//Timer digit 10,000's
	case((timer/10000)%10)
	0:
		begin
		mem[0][105][4:0] = 5'b01110;
		mem[0][104][4:0] = 5'b10001;
		mem[0][103][4:0] = 5'b10001;
		mem[0][102][4:0] = 5'b01110;
		end
	1:
		begin
		mem[0][105][4:0] = 5'b10000;
		mem[0][104][4:0] = 5'b11111;
		mem[0][103][4:0] = 5'b10010;
		mem[0][102][4:0] = 5'b00000;
		end
	2:
		begin
		mem[0][105][4:0] = 5'b10010;
		mem[0][104][4:0] = 5'b10101;
		mem[0][103][4:0] = 5'b11001;
		mem[0][102][4:0] = 5'b10010;
		end
	3:
		begin
		mem[0][105][4:0] = 5'b01010;
		mem[0][104][4:0] = 5'b10101;
		mem[0][103][4:0] = 5'b10101;
		mem[0][102][4:0] = 5'b10001;		
		end
	4:
	begin
		mem[0][105][4:0] = 5'b11111;
		mem[0][104][4:0] = 5'b01010;
		mem[0][103][4:0] = 5'b01100;
		mem[0][102][4:0] = 5'b01000;	
	end
	5:
	begin
		mem[0][105][4:0] = 5'b01001;
		mem[0][104][4:0] = 5'b10101;
		mem[0][103][4:0] = 5'b10101;
		mem[0][102][4:0] = 5'b10111;
	end
	6:
	begin
		mem[0][105][4:0] = 5'b01000;
		mem[0][104][4:0] = 5'b10101;
		mem[0][103][4:0] = 5'b10101;
		mem[0][102][4:0] = 5'b01110;
	end
	7:
	begin
		mem[0][105][4:0] = 5'b00011;
		mem[0][104][4:0] = 5'b00101;
		mem[0][103][4:0] = 5'b01001;
		mem[0][102][4:0] = 5'b10001;
	end
	
	8:
	begin
		mem[0][105][4:0] = 5'b01010;
		mem[0][104][4:0] = 5'b10101;
		mem[0][103][4:0] = 5'b10101;
		mem[0][102][4:0] = 5'b01010;
	end
	9: begin
		mem[0][105][4:0] = 5'b01110;
		mem[0][104][4:0] = 5'b10101;
		mem[0][103][4:0] = 5'b10101;
		mem[0][102][4:0] = 5'b00010;
		end
	default : 
		begin
		mem[0][105][4:0] = 5'b01110;
		mem[0][104][4:0] = 5'b10001;
		mem[0][103][4:0] = 5'b10001;
		mem[0][102][4:0] = 5'b01110;
	end
	endcase
	
	
	//Timer digit 1000's
	case((timer/1000)%10)
	0:
		begin
		mem[0][110][4:0] = 5'b01110;
		mem[0][109][4:0] = 5'b10001;
		mem[0][108][4:0] = 5'b10001;
		mem[0][107][4:0] = 5'b01110;
		end
	1:
		begin
		mem[0][110][4:0] = 5'b10000;
		mem[0][109][4:0] = 5'b11111;
		mem[0][108][4:0] = 5'b10010;
		mem[0][107][4:0] = 5'b00000;
		end
	2:
		begin
		mem[0][110][4:0] = 5'b10010;
		mem[0][109][4:0] = 5'b10101;
		mem[0][108][4:0] = 5'b11001;
		mem[0][107][4:0] = 5'b10010;
		end
	3:
		begin
		mem[0][110][4:0] = 5'b01010;
		mem[0][109][4:0] = 5'b10101;
		mem[0][108][4:0] = 5'b10101;
		mem[0][107][4:0] = 5'b10001;		
		end
	4:
	begin
		mem[0][110][4:0] = 5'b11111;
		mem[0][109][4:0] = 5'b01010;
		mem[0][108][4:0] = 5'b01100;
		mem[0][107][4:0] = 5'b01000;	
	end
	5:
	begin
		mem[0][110][4:0] = 5'b01001;
		mem[0][109][4:0] = 5'b10101;
		mem[0][108][4:0] = 5'b10101;
		mem[0][107][4:0] = 5'b10111;
	end
	6:
	begin
		mem[0][110][4:0] = 5'b01000;
		mem[0][109][4:0] = 5'b10101;
		mem[0][108][4:0] = 5'b10101;
		mem[0][107][4:0] = 5'b01110;
	end
	7:
	begin
		mem[0][110][4:0] = 5'b00011;
		mem[0][109][4:0] = 5'b00101;
		mem[0][108][4:0] = 5'b01001;
		mem[0][107][4:0] = 5'b10001;
	end
	
	8:
	begin
		mem[0][110][4:0] = 5'b01010;
		mem[0][109][4:0] = 5'b10101;
		mem[0][108][4:0] = 5'b10101;
		mem[0][107][4:0] = 5'b01010;
	end
	9: begin
		mem[0][110][4:0] = 5'b01110;
		mem[0][109][4:0] = 5'b10101;
		mem[0][108][4:0] = 5'b10101;
		mem[0][107][4:0] = 5'b00010;
		end
	default : 
		begin
		mem[0][110][4:0] = 5'b01110;
		mem[0][109][4:0] = 5'b10001;
		mem[0][108][4:0] = 5'b10001;
		mem[0][107][4:0] = 5'b01110;
	end
	endcase
	
	
	//Timer digit 100's
	case((timer/100)%10)
	0:
		begin
		mem[0][115][4:0] = 5'b01110;
		mem[0][114][4:0] = 5'b10001;
		mem[0][113][4:0] = 5'b10001;
		mem[0][112][4:0] = 5'b01110;
		end
	1:
		begin
		mem[0][115][4:0] = 5'b10000;
		mem[0][114][4:0] = 5'b11111;
		mem[0][113][4:0] = 5'b10010;
		mem[0][112][4:0] = 5'b00000;
		end
	2:
		begin
		mem[0][115][4:0] = 5'b10010;
		mem[0][114][4:0] = 5'b10101;
		mem[0][113][4:0] = 5'b11001;
		mem[0][112][4:0] = 5'b10010;
		end
	3:
		begin
		mem[0][115][4:0] = 5'b01010;
		mem[0][114][4:0] = 5'b10101;
		mem[0][113][4:0] = 5'b10101;
		mem[0][112][4:0] = 5'b10001;		
		end
	4:
	begin
		mem[0][115][4:0] = 5'b11111;
		mem[0][114][4:0] = 5'b01010;
		mem[0][113][4:0] = 5'b01100;
		mem[0][112][4:0] = 5'b01000;	
	end
	5:
	begin
		mem[0][115][4:0] = 5'b01001;
		mem[0][114][4:0] = 5'b10101;
		mem[0][113][4:0] = 5'b10101;
		mem[0][112][4:0] = 5'b10111;
	end
	6:
	begin
		mem[0][115][4:0] = 5'b01000;
		mem[0][114][4:0] = 5'b10101;
		mem[0][113][4:0] = 5'b10101;
		mem[0][112][4:0] = 5'b01110;
	end
	7:
	begin
		mem[0][115][4:0] = 5'b00011;
		mem[0][114][4:0] = 5'b00101;
		mem[0][113][4:0] = 5'b01001;
		mem[0][112][4:0] = 5'b10001;
	end
	
	8:
	begin
		mem[0][115][4:0] = 5'b01010;
		mem[0][114][4:0] = 5'b10101;
		mem[0][113][4:0] = 5'b10101;
		mem[0][112][4:0] = 5'b01010;
	end
	9: begin
		mem[0][115][4:0] = 5'b01110;
		mem[0][114][4:0] = 5'b10101;
		mem[0][113][4:0] = 5'b10101;
		mem[0][112][4:0] = 5'b00010;
		end
	default : 
		begin
		mem[0][115][4:0] = 5'b01110;
		mem[0][114][4:0] = 5'b10001;
		mem[0][113][4:0] = 5'b10001;
		mem[0][112][4:0] = 5'b01110;
	end
	endcase
	
	
	//Timer digit 10's
	case((timer/10)%10)
	0:
		begin
		mem[0][120][4:0] = 5'b01110;
		mem[0][119][4:0] = 5'b10001;
		mem[0][118][4:0] = 5'b10001;
		mem[0][117][4:0] = 5'b01110;
		end
	1:
		begin
		mem[0][120][4:0] = 5'b10000;
		mem[0][119][4:0] = 5'b11111;
		mem[0][118][4:0] = 5'b10010;
		mem[0][117][4:0] = 5'b00000;
		end
	2:
		begin
		mem[0][120][4:0] = 5'b10010;
		mem[0][119][4:0] = 5'b10101;
		mem[0][118][4:0] = 5'b11001;
		mem[0][117][4:0] = 5'b10010;
		end
	3:
		begin
		mem[0][120][4:0] = 5'b01010;
		mem[0][119][4:0] = 5'b10101;
		mem[0][118][4:0] = 5'b10101;
		mem[0][117][4:0] = 5'b10001;		
		end
	4:
	begin
		mem[0][120][4:0] = 5'b11111;
		mem[0][119][4:0] = 5'b01010;
		mem[0][118][4:0] = 5'b01100;
		mem[0][117][4:0] = 5'b01000;	
	end
	5:
	begin
		mem[0][120][4:0] = 5'b01001;
		mem[0][119][4:0] = 5'b10101;
		mem[0][118][4:0] = 5'b10101;
		mem[0][117][4:0] = 5'b10111;
	end
	6:
	begin
		mem[0][120][4:0] = 5'b01000;
		mem[0][119][4:0] = 5'b10101;
		mem[0][118][4:0] = 5'b10101;
		mem[0][117][4:0] = 5'b01110;
	end
	7:
	begin
		mem[0][120][4:0] = 5'b00011;
		mem[0][119][4:0] = 5'b00101;
		mem[0][118][4:0] = 5'b01001;
		mem[0][117][4:0] = 5'b10001;
	end
	
	8:
	begin
		mem[0][120][4:0] = 5'b01010;
		mem[0][119][4:0] = 5'b10101;
		mem[0][118][4:0] = 5'b10101;
		mem[0][117][4:0] = 5'b01010;
	end
	9: begin
		mem[0][120][4:0] = 5'b01110;
		mem[0][119][4:0] = 5'b10101;
		mem[0][118][4:0] = 5'b10101;
		mem[0][117][4:0] = 5'b00010;
		end
	default : 
		begin
		mem[0][120][4:0] = 5'b01110;
		mem[0][119][4:0] = 5'b10001;
		mem[0][118][4:0] = 5'b10001;
		mem[0][117][4:0] = 5'b01110;
	end
	endcase
	
	//Timer digit 1's
	case(timer%10)
	0:
		begin
		mem[0][125][4:0] = 5'b01110;
		mem[0][124][4:0] = 5'b10001;
		mem[0][123][4:0] = 5'b10001;
		mem[0][122][4:0] = 5'b01110;
		end
	1:
		begin
		mem[0][125][4:0] = 5'b10000;
		mem[0][124][4:0] = 5'b11111;
		mem[0][123][4:0] = 5'b10010;
		mem[0][122][4:0] = 5'b00000;
		end
	2:
		begin
		mem[0][125][4:0] = 5'b10010;
		mem[0][124][4:0] = 5'b10101;
		mem[0][123][4:0] = 5'b11001;
		mem[0][122][4:0] = 5'b10010;
		end
	3:
		begin
		mem[0][125][4:0] = 5'b01010;
		mem[0][124][4:0] = 5'b10101;
		mem[0][123][4:0] = 5'b10101;
		mem[0][122][4:0] = 5'b10001;		
		end
	4:
	begin
		mem[0][125][4:0] = 5'b11111;
		mem[0][124][4:0] = 5'b01010;
		mem[0][123][4:0] = 5'b01100;
		mem[0][122][4:0] = 5'b01000;	
	end
	5:
	begin
		mem[0][125][4:0] = 5'b01001;
		mem[0][124][4:0] = 5'b10101;
		mem[0][123][4:0] = 5'b10101;
		mem[0][122][4:0] = 5'b10111;
	end
	6:
	begin
		mem[0][125][4:0] = 5'b01000;
		mem[0][124][4:0] = 5'b10101;
		mem[0][123][4:0] = 5'b10101;
		mem[0][122][4:0] = 5'b01110;
	end
	7:
	begin
		mem[0][125][4:0] = 5'b00011;
		mem[0][124][4:0] = 5'b00101;
		mem[0][123][4:0] = 5'b01001;
		mem[0][122][4:0] = 5'b10001;
	end
	
	8:
	begin
		mem[0][125][4:0] = 5'b01010;
		mem[0][124][4:0] = 5'b10101;
		mem[0][123][4:0] = 5'b10101;
		mem[0][122][4:0] = 5'b01010;
	end
	9: begin
		mem[0][125][4:0] = 5'b01110;
		mem[0][124][4:0] = 5'b10101;
		mem[0][123][4:0] = 5'b10101;
		mem[0][122][4:0] = 5'b00010;
		end
	default : 
		begin
		mem[0][125][4:0] = 5'b01110;
		mem[0][124][4:0] = 5'b10001;
		mem[0][123][4:0] = 5'b10001;
		mem[0][122][4:0] = 5'b01110;
	end
	endcase
	end		
	end
//First lane Divider 20
	always@(negedge clk_1) begin
	if (init1 == 0) begin
		
/*		mem[1][0] = 8'b00110000;
		mem[1][1] = 8'b11111100;
		mem[1][2] = 8'b11111100;
		mem[1][3] = 8'b00110000;
		mem[1][4] = 8'b11111100;
		mem[1][5] = 8'b11001100;
*/		
		mem[1][15] = 8'b00110000;
		mem[1][16] = 8'b11111100;
		mem[1][17] = 8'b11111100;
		mem[1][18] = 8'b00110000;
		mem[1][19] = 8'b11111100;
		mem[1][20] = 8'b11001100;

/*		
		mem[1][50] = 8'b00110000;
		mem[1][51] = 8'b11111100;
		mem[1][52] = 8'b11111100;
		mem[1][53] = 8'b00110000;
		mem[1][54] = 8'b11111100;
		mem[1][55] = 8'b11001100;
*/		
		mem[1][70] = 8'b00110000;
		mem[1][71] = 8'b11111100;
		mem[1][72] = 8'b11111100;
		mem[1][73] = 8'b00110000;
		mem[1][74] = 8'b11111100;
		mem[1][75] = 8'b11001100;
		
		mem[1][140] = 8'b00110000;
		mem[1][141] = 8'b11111100;
		mem[1][142] = 8'b11111100;
		mem[1][143] = 8'b00110000;
		mem[1][144] = 8'b11111100;
		mem[1][145] = 8'b11001100;

/*		mem[1][188] = 8'b00110000;
		mem[1][189] = 8'b11111100;
		mem[1][190] = 8'b11111100;
		mem[1][191] = 8'b00110000;
		mem[1][192] = 8'b11111100;
		mem[1][193] = 8'b11001100;
*/		
		mem[1][225] = 8'b00110000;
		mem[1][226] = 8'b11111100;
		mem[1][227] = 8'b11111100;
		mem[1][228] = 8'b00110000;
		mem[1][229] = 8'b11111100;
		mem[1][230] = 8'b11001100;
				
		init1 = 1;
	end
		temp1[7:0] = mem[1][0][7:0] ;
		for ( move1 = 0; move1 < 255 ; move1 = move1+1) begin
			mem[1][move1][7:0] = mem[1][move1+1][7:0] ;
		end
		mem[1][255][7:0] = temp1[7:0];
end
//Second Lane 21
	always@(negedge clk_2) begin
	if (init2 == 0) begin
/*		mem[2][0] = 8'b00110000;
		mem[2][1] = 8'b11111100;
		mem[2][2] = 8'b11111100;
		mem[2][3] = 8'b00110000;
		mem[2][4] = 8'b11111100;
		mem[2][5] = 8'b11001100;
*/		
		mem[2][17] = 8'b00110000;
		mem[2][18] = 8'b11111100;
		mem[2][19] = 8'b11111100;
		mem[2][20] = 8'b00110000;
		mem[2][21] = 8'b11111100;
		mem[2][22] = 8'b11001100;
/*	
		mem[2][32] = 8'b00110000;
		mem[2][33] = 8'b11111100;
		mem[2][34] = 8'b11111100;
		mem[2][35] = 8'b00110000;
		mem[2][36] = 8'b11111100;
		mem[2][37] = 8'b11001100;
		
		mem[2][46] = 8'b00110000;
		mem[2][47] = 8'b11111100;
		mem[2][48] = 8'b11111100;
		mem[2][49] = 8'b00110000;
		mem[2][50] = 8'b11111100;
		mem[2][51] = 8'b11001100;
		
		mem[2][75] = 8'b00110000;
		mem[2][76] = 8'b11111100;
		mem[2][77] = 8'b11111100;
		mem[2][78] = 8'b00110000;
		mem[2][79] = 8'b11111100;
		mem[2][80] = 8'b11001100;
*/				
		mem[2][111] = 8'b00110000;
		mem[2][112] = 8'b11111100;
		mem[2][113] = 8'b11111100;
		mem[2][114] = 8'b00110000;
		mem[2][115] = 8'b11111100;
		mem[2][116] = 8'b11001100;
		
		mem[2][175] = 8'b00110000;
		mem[2][176] = 8'b11111100;
		mem[2][177] = 8'b11111100;
		mem[2][178] = 8'b00110000;
		mem[2][179] = 8'b11111100;
		mem[2][180] = 8'b11001100;
						
		init2 = 1;
	end
		temp2[7:0] = mem[2][0][7:0] ;
		for ( move2 = 0; move2 < 255 ; move2 = move2+1) begin
			mem[2][move2][7:0] = mem[2][move2+1][7:0] ;
		end
		mem[2][255][7:0] = temp2[7:0];
end
//Third lane  22
	always@(negedge clk_3) begin
	if (init3 == 0) begin
/*		mem[3][0] = 8'b00110000;
		mem[3][1] = 8'b11111100;
		mem[3][2] = 8'b11111100;
		mem[3][3] = 8'b00110000;
		mem[3][4] = 8'b11111100;
		mem[3][5] = 8'b11001100;
		
		mem[3][25] = 8'b00110000;
		mem[3][26] = 8'b11111100;
		mem[3][27] = 8'b11111100;
		mem[3][28] = 8'b00110000;
		mem[3][29] = 8'b11111100;
		mem[3][30] = 8'b11001100;
*/		
		mem[3][55] = 8'b00110000;
		mem[3][56] = 8'b11111100;
		mem[3][57] = 8'b11111100;
		mem[3][58] = 8'b00110000;
		mem[3][59] = 8'b11111100;
		mem[3][60] = 8'b11001100;
		
		mem[3][80] = 8'b00110000;
		mem[3][81] = 8'b11111100;
		mem[3][82] = 8'b11111100;
		mem[3][83] = 8'b00110000;
		mem[3][84] = 8'b11111100;
		mem[3][85] = 8'b11001100;
		
		mem[3][168] = 8'b00110000;
		mem[3][169] = 8'b11111100;
		mem[3][170] = 8'b11111100;
		mem[3][171] = 8'b00110000;
		mem[3][172] = 8'b11111100;
		mem[3][173] = 8'b11001100;
		
		mem[3][211] = 8'b00110000;
		mem[3][212] = 8'b11111100;
		mem[3][213] = 8'b11111100;
		mem[3][214] = 8'b00110000;
		mem[3][215] = 8'b11111100;
		mem[3][216]= 8'b11001100;
				
		init3 = 1;
	end
		temp3[7:0] = mem[3][0][7:0] ;
		for ( move3 = 0; move3 < 255 ; move3 = move3+1) begin
			mem[3][move3][7:0] = mem[3][move3+1][7:0] ;
		end
		mem[3][255][7:0] = temp3[7:0];
end
//Fourth lane 21
	always@(negedge clk_4) begin
	if (init4 == 0) begin
		mem[4][0] = 8'b00110000;
		mem[4][1] = 8'b11111100;
		mem[4][2] = 8'b11111100;
		mem[4][3] = 8'b00110000;
		mem[4][4] = 8'b11111100;
		mem[4][5] = 8'b11001100;
		
/*		mem[4][45] = 8'b00110000;
		mem[4][46] = 8'b11111100;
		mem[4][47] = 8'b11111100;
		mem[4][48] = 8'b00110000;
		mem[4][49] = 8'b11111100;
		mem[4][50] = 8'b11001100;
		
		mem[4][65] = 8'b00110000;
		mem[4][66] = 8'b11111100;
		mem[4][67] = 8'b11111100;
		mem[4][68] = 8'b00110000;
		mem[4][69] = 8'b11111100;
		mem[4][70] = 8'b11001100;
*/		
		mem[4][115] = 8'b00110000;
		mem[4][116] = 8'b11111100;
		mem[4][117] = 8'b11111100;
		mem[4][118] = 8'b00110000;
		mem[4][119] = 8'b11111100;
		mem[4][120] = 8'b11001100;
		
		mem[4][145] = 8'b00110000;
		mem[4][146] = 8'b11111100;
		mem[4][147] = 8'b11111100;
		mem[4][148] = 8'b00110000;
		mem[4][149] = 8'b11111100;
		mem[4][150] = 8'b11001100;
		
		mem[4][200] = 8'b00110000;
		mem[4][201] = 8'b11111100;
		mem[4][202] = 8'b11111100;
		mem[4][203] = 8'b00110000;
		mem[4][204] = 8'b11111100;
		mem[4][205] = 8'b11001100;
		
		mem[4][237] = 8'b00110000;
		mem[4][238] = 8'b11111100;
		mem[4][239] = 8'b11111100;
		mem[4][240] = 8'b00110000;
		mem[4][241] = 8'b11111100;
		mem[4][242] = 8'b11001100;
		
		
		init4 = 1;
	end
		temp4[7:0] = mem[4][0][7:0] ;
		for ( move4 = 0; move4 < 255 ; move4 = move4+1) begin
			mem[4][move4][7:0] = mem[4][move4+1][7:0] ;
		end
		mem[4][255][7:0] = temp4[7:0];
	
end
//Fifth lane 23
	always@(negedge clk_5) begin
	if (init5 == 0) begin
/*		mem[5][21] = 8'b00110000;
		mem[5][22] = 8'b11111100;
		mem[5][23] = 8'b11111100;
		mem[5][24] = 8'b00110000;
		mem[5][25] = 8'b11111100;
		mem[5][26] = 8'b11001100;
*/		
		mem[5][33] = 8'b00110000;
		mem[5][34] = 8'b11111100;
		mem[5][35] = 8'b11111100;
		mem[5][37] = 8'b00110000;
		mem[5][38] = 8'b11111100;
		mem[5][39] = 8'b11001100;
		
/*		
		mem[5][45] = 8'b00110000;
		mem[5][46] = 8'b11111100;
		mem[5][47] = 8'b11111100;
		mem[5][48] = 8'b00110000;
		mem[5][49] = 8'b11111100;
		mem[5][50] = 8'b11001100;
*/	
		mem[5][58] = 8'b00110000;
		mem[5][59] = 8'b11111100;
		mem[5][60] = 8'b11111100;
		mem[5][61] = 8'b00110000;
		mem[5][62] = 8'b11111100;
		mem[5][63] = 8'b11001100;
		
		mem[5][75] = 8'b00110000;
		mem[5][76] = 8'b11111100;
		mem[5][77] = 8'b11111100;
		mem[5][78] = 8'b00110000;
		mem[5][79] = 8'b11111100;
		mem[5][80] = 8'b11001100;
/*
		mem[5][100] = 8'b00110000;
		mem[5][101] = 8'b11111100;
		mem[5][102] = 8'b11111100;
		mem[5][103] = 8'b00110000;
		mem[5][104] = 8'b11111100;
		mem[5][105] = 8'b11001100;
/*	
		mem[5][115] = 8'b00110000;
		mem[5][116] = 8'b11111100;
		mem[5][117] = 8'b11111100;
		mem[5][118] = 8'b00110000;
		mem[5][119] = 8'b11111100;
		mem[5][120] = 8'b11001100;
*/		
		mem[5][130] = 8'b00110000;
		mem[5][131] = 8'b11111100;
		mem[5][132] = 8'b11111100;
		mem[5][133] = 8'b00110000;
		mem[5][134] = 8'b11111100;
		mem[5][135] = 8'b11001100;
		
/*		mem[5][160] = 8'b00110000;
		mem[5][161] = 8'b11111100;
		mem[5][162] = 8'b11111100;
		mem[5][163] = 8'b00110000;
		mem[5][164] = 8'b11111100;
		mem[5][165] = 8'b11001100;
*/		
		mem[5][182] = 8'b00110000;
		mem[5][183] = 8'b11111100;
		mem[5][184] = 8'b11111100;
		mem[5][185] = 8'b00110000;
		mem[5][186] = 8'b11111100;
		mem[5][187] = 8'b11001100;
		
/*		mem[5][199] = 8'b00110000;
		mem[5][200] = 8'b11111100;
		mem[5][201] = 8'b11111100;
		mem[5][202] = 8'b00110000;
		mem[5][203] = 8'b11111100;
		mem[5][204] = 8'b11001100;
		
		mem[5][220] = 8'b00110000;
		mem[5][221] = 8'b11111100;
		mem[5][222] = 8'b11111100;
		mem[5][223] = 8'b00110000;
		mem[5][224] = 8'b11111100;
		mem[5][225] = 8'b11001100;
/*		
		mem[5][245] = 8'b00110000;
		mem[5][246] = 8'b11111100;
		mem[5][247] = 8'b11111100;
		mem[5][248] = 8'b00110000;
		mem[5][249] = 8'b11111100;
		mem[5][250] = 8'b11001100;
*/		
		init5 = 1;
	end
		temp5[7:0] = mem[5][0][7:0] ;
		for ( move5 = 0; move5 < 255 ; move5 = move5+1) begin
			mem[5][move5][7:0] = mem[5][move5+1][7:0] ;
		end
		mem[5][255][7:0] = temp5[7:0];
	
end
//Sixth lane 20
	always@(negedge clk_6) begin
	if (init6 == 0) begin
		mem[6][10] = 8'b00110000;
		mem[6][11] = 8'b11111100;
		mem[6][12] = 8'b11111100;
		mem[6][13] = 8'b00110000;
		mem[6][14] = 8'b11111100;
		mem[6][15] = 8'b11001100;
/*		
		mem[6][35] = 8'b00110000;
		mem[6][36] = 8'b11111100;
		mem[6][37] = 8'b11111100;
		mem[6][38] = 8'b00110000;
		mem[6][39] = 8'b11111100;
		mem[6][40] = 8'b11001100;
*/		
		mem[6][60] = 8'b00110000;
		mem[6][61] = 8'b11111100;
		mem[6][62] = 8'b11111100;
		mem[6][63] = 8'b00110000;
		mem[6][64] = 8'b11111100;
		mem[6][65] = 8'b11001100;
/*		
		mem[6][110] = 8'b00110000;
		mem[6][111] = 8'b11111100;
		mem[6][112] = 8'b11111100;
		mem[6][113] = 8'b00110000;
		mem[6][114] = 8'b11111100;
		mem[6][115] = 8'b11001100;
		
		mem[6][133] = 8'b00110000;
		mem[6][134] = 8'b11111100;
		mem[6][135] = 8'b11111100;
		mem[6][136] = 8'b00110000;
		mem[6][137] = 8'b11111100;
		mem[6][138] = 8'b11001100;
		
		mem[6][170] = 8'b00110000;
		mem[6][171] = 8'b11111100;
		mem[6][172] = 8'b11111100;
		mem[6][173] = 8'b00110000;
		mem[6][174] = 8'b11111100;
		mem[6][175] = 8'b11001100;
		
*/		
		mem[6][200] = 8'b00110000;
		mem[6][201] = 8'b11111100;
		mem[6][202] = 8'b11111100;
		mem[6][203] = 8'b00110000;
		mem[6][204] = 8'b11111100;
		mem[6][205] = 8'b11001100;
		
		
		init6 = 1;
	end
		temp6[7:0] = mem[6][0][7:0] ;
		for ( move6 = 0; move6 < 255; move6 = move6+1) begin
			mem[6][move6][7:0] = mem[6][move6+1][7:0] ;
		end
		mem[6][255][7:0] = temp6[7:0];
		
end
//Seventh lane 22
	always@(negedge clk_7) begin
	if (init7 == 0) begin
/*		mem[7][1] = 8'b00110000;
		mem[7][2] = 8'b11111100;
		mem[7][3] = 8'b11111100;
		mem[7][4] = 8'b00110000;
		mem[7][5] = 8'b11111100;
		mem[7][7] = 8'b11001100;
			
		mem[7][15] = 8'b00110000;
		mem[7][16] = 8'b11111100;
		mem[7][17] = 8'b11111100;
		mem[7][18] = 8'b00110000;
		mem[7][19] = 8'b11111100;
		mem[7][20] = 8'b11001100;
		
*/
		mem[7][25] = 8'b00110000;
		mem[7][26] = 8'b11111100;
		mem[7][27] = 8'b11111100;
		mem[7][28] = 8'b00110000;
		mem[7][29] = 8'b11111100;
		mem[7][30] = 8'b11001100;
/*		
		mem[7][60] = 8'b00110000;
		mem[7][61] = 8'b11111100;
		mem[7][62] = 8'b11111100;
		mem[7][63] = 8'b00110000;
		mem[7][64] = 8'b11111100;
		mem[7][65] = 8'b11001100;
*/		
		mem[7][91] = 8'b00110000;
		mem[7][92] = 8'b11111100;
		mem[7][93] = 8'b11111100;
		mem[7][94] = 8'b00110000;
		mem[7][95] = 8'b11111100;
		mem[7][96] = 8'b11001100;
/*		
		mem[7][135] = 8'b00110000;
		mem[7][136] = 8'b11111100;
		mem[7][137] = 8'b11111100;
		mem[7][138] = 8'b00110000;
		mem[7][139] = 8'b11111100;
		mem[7][140] = 8'b11001100;
*/		
		mem[7][150] = 8'b00110000;
		mem[7][151] = 8'b11111100;
		mem[7][152] = 8'b11111100;
		mem[7][153] = 8'b00110000;
		mem[7][154] = 8'b11111100;
		mem[7][155] = 8'b11001100;
		
/*		mem[7][190] = 8'b00110000;
		mem[7][191] = 8'b11111100;
		mem[7][192] = 8'b11111100;
		mem[7][193] = 8'b00110000;
		mem[7][194] = 8'b11111100;
		mem[7][195] = 8'b11001100;
		
/*		mem[7][225] = 8'b00110000;
		mem[7][226] = 8'b11111100;
		mem[7][227] = 8'b11111100;
		mem[7][228] = 8'b00110000;
		mem[7][229] = 8'b11111100;
		mem[7][230] = 8'b11001100;
*/		
		init7 = 1;
	end
		temp7[7:0] = mem[7][0][7:0] ;
		for ( move7 = 0; move7 < 255 ; move7 = move7+1) begin
			mem[7][move7][7:0] = mem[7][move7+1][7:0] ;
		end
		mem[7][255][7:0] = temp7[7:0];
		
end
//Clock dividing function
always @ (posedge clk) divider <= divider + 1;
//Screen Refreshing block
always@(posedge divider[8]) begin
		count <= count + 1;
		reset <= 1;
		//cs1 <= 1; 
		//cs2 <= 1;
		
		if(count <= 9)
			begin cs1<=1; cs2<=1;lcd_rs <= 0; lcd_rw <= 0; lcd_e <= 0; lcd_data <= 8'b00000000; end
		else if(count == 10)
			begin lcd_rs <= 0; lcd_rw <= 0; lcd_data <= 8'b00111111; lcd_e <= 1; end
		else if(count == 11)
			lcd_e <= 0;
		else if(count == 12)
			begin cs1<=1;cs2<=1;lcd_rs <= 0; lcd_rw <= 0; lcd_data <= 184+page; lcd_e <= 1; end
		else if(count == 13)
			lcd_e <= 0;
		else if(count == 14)
			begin lcd_rs <= 0; lcd_rw <= 0; lcd_data <= 64+col ; lcd_e <= 1; end
		else if(count == 15)
			lcd_e <= 0;
		else begin		
			if(!already_on) begin
				if(gameover==0 && start==0 )begin 
				if (i <64 ) begin
					cs1 <= 1;
					cs2 <= 0;
				end 
				else if (i > 63) begin
					cs1 <= 0;
					cs2 <= 1;
				end
				
				lcd_rs <=1 ; 
				lcd_rw <= 0; 
				if (i<6) begin 
					if((carmem[page][i]>0)&& (mem[page][i]>0))
						gameover = 1 ; 
					else lcd_data = carmem[page][i] | mem [page][i] ; 
				end
				if (i>=6 && i<128) begin  lcd_data = mem[page][i] ; end 
				lcd_e <= 1; 
				i <= i+1;
				already_on <= 1;
				if (i == 128) begin
					i <= 0;
					page = (page ==7)? 0 : page+ 1 ;
					count <= 10;
				end
				end
				else if((gameover==1 ) | (start == 1)) begin 
				if (i <64 ) begin
					cs1 <= 1;
					cs2 <= 0;
				end 
				else if (i > 63) begin
					cs1 <= 0;
					cs2 <= 1;
				end
				
				lcd_rs <=1 ; 
				lcd_rw <= 0; 
				lcd_data = tmem[page][i];
				lcd_e <= 1; 
				i <= i+1;
				already_on <= 1;
				if (i == 128) begin
					i <= 0;
					page = (page ==7)? 0 : page+ 1 ;
					count <= 10;
				end
				end
			end
			else begin
				already_on <= 0;
				lcd_e <= 0;
			end
		end
end		

//Welcome and Game Over 
always@(negedge divider[21]) begin
	if((timer1<50) && (init_w==0) && (init_g==1)) begin 
	//Letter W
	tmem[3][43][4:0] = 5'b11111; 
	tmem[3][44][4:0] = 5'b10000; 
	tmem[3][45][4:0] = 5'b11100; 
	tmem[3][46][4:0] = 5'b10000; 
	tmem[3][47][4:0] = 5'b11111;

//Letter E 
	tmem[3][49][4:0] = 5'b11111; 
	tmem[3][50][4:0] = 5'b10101; 
	tmem[3][51][4:0] = 5'b10101;
	tmem[3][52][4:0] = 5'b10101;
	tmem[3][53][4:0] = 5'b10001;
	
//Letter L	
	tmem[3][55][4:0] = 5'b11111; 
	tmem[3][56][4:0] = 5'b10000; 
	tmem[3][57][4:0] = 5'b10000; 
	tmem[3][58][4:0] = 5'b10000; 
	tmem[3][59][4:0] = 5'b10000;

//Letter "C"
	tmem[3][61][4:0] = 5'b00100; 
	tmem[3][62][4:0] = 5'b01010; 
	tmem[3][63][4:0] = 5'b10001;
	tmem[3][64][4:0] = 5'b10001;
	tmem[3][65][4:0] = 5'b10001;	

//Letter "O"
	tmem[3][67][4:0] = 5'b01110; 
	tmem[3][68][4:0] = 5'b10001; 
	tmem[3][69][4:0] = 5'b10001;
	tmem[3][70][4:0] = 5'b10001;
	tmem[3][71][4:0] = 5'b01110;
	
//Letter M
	tmem[3][73][4:0] = 5'b11111; 
	tmem[3][74][4:0] = 5'b00010; 
	tmem[3][75][4:0] = 5'b00100; 
	tmem[3][76][4:0] = 5'b00010; 
	tmem[3][77][4:0] = 5'b11111;
	
//Letter E 
	tmem[3][79][4:0] = 5'b11111; 
	tmem[3][80][4:0] = 5'b10101; 
	tmem[3][81][4:0] = 5'b10101;
	tmem[3][82][4:0] = 5'b10101;
	tmem[3][83][4:0] = 5'b10001;

//Letter T 
	tmem[4][55][4:0] = 5'b00001; 
	tmem[4][56][4:0] = 5'b00001; 
	tmem[4][57][4:0] = 5'b11111;
	tmem[4][58][4:0] = 5'b00001;
	tmem[4][59][4:0] = 5'b00001;

//Letter "O"
	tmem[4][61][4:0] = 5'b01110; 
	tmem[4][62][4:0] = 5'b10001; 
	tmem[4][63][4:0] = 5'b10001;
	tmem[4][64][4:0] = 5'b10001;
	tmem[4][65][4:0] = 5'b01110;
	
//Letter "C"
	tmem[5][40][4:0] = 5'b00100; 
	tmem[5][41][4:0] = 5'b01010; 
	tmem[5][42][4:0] = 5'b10001;
	tmem[5][43][4:0] = 5'b10001;
	tmem[5][44][4:0] = 5'b10001;	
	
//Letter A
	tmem[5][46][4:0] = 5'b11110; 
	tmem[5][47][4:0] = 5'b00101; 
	tmem[5][48][4:0] = 5'b00101; 
	tmem[5][49][4:0] = 5'b00101; 
	tmem[5][50][4:0] = 5'b11110;	

//Letter R 	
	tmem[5][52][4:0] = 5'b11111; 
	tmem[5][53][4:0] = 5'b00101; 
	tmem[5][54][4:0] = 5'b00101;
	tmem[5][55][4:0] = 5'b01010;
	tmem[5][56][4:0] = 5'b10000;
	
//Letter G
	tmem[5][61][4:0] = 5'b11111; 
	tmem[5][62][4:0] = 5'b10001; 
	tmem[5][63][4:0] = 5'b10001; 
	tmem[5][64][4:0] = 5'b10101; 
	tmem[5][65][4:0] = 5'b11101;
	
//Letter A
	tmem[5][67][4:0] = 5'b11110; 
	tmem[5][68][4:0] = 5'b00101; 
	tmem[5][69][4:0] = 5'b00101; 
	tmem[5][70][4:0] = 5'b00101; 
	tmem[5][71][4:0] = 5'b11110;
	
//Letter M
	tmem[5][73][4:0] = 5'b11111; 
	tmem[5][74][4:0] = 5'b00010; 
	tmem[5][75][4:0] = 5'b00100; 
	tmem[5][76][4:0] = 5'b00010; 
	tmem[5][77][4:0] = 5'b11111;

//Letter E 
	tmem[5][79][4:0] = 5'b11111; 
	tmem[5][80][4:0] = 5'b10101; 
	tmem[5][81][4:0] = 5'b10101;
	tmem[5][82][4:0] = 5'b10101;
	tmem[5][83][4:0] = 5'b10001;	
	
	end
	else if ((timer1 >=50) && (init_w==0) && (init_g==1)) init_w = 1; 
	else if((timer1 >=50)&& (init_g==1) && (init_w==1)) begin for (i1=3; i1<=5; i1=i1+1)begin for(j1=0; j1<=127; j1=j1+1) begin tmem[i1][j1][4:0]=5'b00000; end end init_g=0; end 
	else if((timer1 >=50) && (init_g==0) && (gameover==0)) begin 
		
//Letter G
	tmem[4][41][4:0] = 5'b11111; 
	tmem[4][42][4:0] = 5'b10001; 
	tmem[4][43][4:0] = 5'b10001; 
	tmem[4][44][4:0] = 5'b10101; 
	tmem[4][45][4:0] = 5'b11101;
	
//Letter A
	tmem[4][47][4:0] = 5'b11110; 
	tmem[4][48][4:0] = 5'b00101; 
	tmem[4][49][4:0] = 5'b00101; 
	tmem[4][50][4:0] = 5'b00101; 
	tmem[4][51][4:0] = 5'b11110;
	
//Letter M
	tmem[4][53][4:0] = 5'b11111; 
	tmem[4][54][4:0] = 5'b00010; 
	tmem[4][55][4:0] = 5'b00100; 
	tmem[4][56][4:0] = 5'b00010; 
	tmem[4][57][4:0] = 5'b11111;

//Letter E 
	tmem[4][59][4:0] = 5'b11111; 
	tmem[4][80][4:0] = 5'b10101; 
	tmem[4][61][4:0] = 5'b10101;
	tmem[4][62][4:0] = 5'b10101;
	tmem[4][63][4:0] = 5'b10001;
	
//Letter O
	tmem[4][67][4:0] = 5'b01110; 
	tmem[4][68][4:0] = 5'b10001; 
	tmem[4][69][4:0] = 5'b10001;
	tmem[4][70][4:0] = 5'b10001;
	tmem[4][71][4:0] = 5'b01110;
	
//Letter V 
	tmem[4][73][4:0] = 5'b00011; 
	tmem[4][74][4:0] = 5'b01100; 
	tmem[4][75][4:0] = 5'b10000;
	tmem[4][76][4:0] = 5'b01100;
	tmem[4][77][4:0] = 5'b00011;
	
//Letter E 
	tmem[4][79][4:0] = 5'b11111; 
	tmem[4][80][4:0] = 5'b10101; 
	tmem[4][81][4:0] = 5'b10101;
	tmem[4][82][4:0] = 5'b10101;
	tmem[4][83][4:0] = 5'b10001;

//Letter R 	
	tmem[4][85][4:0] = 5'b11111; 
	tmem[4][86][4:0] = 5'b00101; 
	tmem[4][87][4:0] = 5'b00101;
	tmem[4][88][4:0] = 5'b01010;
	tmem[4][89][4:0] = 5'b10000;

	end
   else if(gameover) begin 
		temp_t[7:0] = tmem[4][0][7:0] ;
		for ( move_t = 0; move_t < 127 ; move_t = move_t+1) begin
			tmem[4][move_t][7:0] = tmem[4][move_t+1][7:0] ;
		end
		tmem[4][127][7:0] = temp_t[7:0];
	end 
end
endmodule
